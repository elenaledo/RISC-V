module decoder (
  input logic clk_i,
  input logic 
);
